// This is header.vh
