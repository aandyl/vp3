`define FOO x22
