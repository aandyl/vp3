module ports (
    input input_scalar,
    input [9:0] input_vector,
    output output_scalar,
    output [9:0] output_vector
);

endmodule
